-- Work in progress
