library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.sha256_pkg.ALL;
use IEEE.NUMERIC_STD.ALL;

entity sha256_core_controller is 
	port(
		clk : in std_logic
		
		
		
		
		
		
		);